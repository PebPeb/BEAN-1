

module top_tb();
  reg clk, reset = 0;

  initial clk <= 0;
	always #1 clk <= ~clk;
	
  top DUT (
    .clk(clk), 
    .reset(reset)
  );

  initial begin
    #200
    $finish;
  end

  integer i;
  initial begin
    $dumpfile("top_tb.vcd");
    $dumpvars(0, top_tb);
    for (i = 0; i < 32; i = i + 1)
      $dumpvars(1, DUT.CPU.data_unit.regFILE.x[i]);
  end
endmodule

